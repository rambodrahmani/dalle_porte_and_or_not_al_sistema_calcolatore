/**
 * File:    RL-20180626.v
 *
 * Author:  Rambod Rahmani <rambodrahmani@autistici.org>
 *          Created on 14/07/2019.
 */

module RL_20180626();
endmodule

