/**
 * File: Riconoscitore_di_Sequenza_Mealy_Ritardato.v
 *       
 * Author: Rambod Rahmani <rambodrahmani@autistici.org>
 *         Created on 12/06/2019.
 */

module Riconoscitore_di_Sequenza_Mealy_Ritardato();
endmodule

